class Packet;

    rand logic [7:0] TX_DATA;

    // Display function.
    


endclass